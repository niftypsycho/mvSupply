C:\DOCUMENTS AND SETTINGS\FFT9ND\DESKTOP\DATA\MY CIRCUITS B\CS5171-2-4\CS5171 (FROM INTUSOFT AND EDITED).CIR SETUP1
*#SAVE V(1) @L2[I] @R7[I] @R7[P] V(FB) @R8[I] @R8[P] @R9[I]
*#SAVE @R9[P] @C3[I] @R10[I] @R10[P] V(11) @C1[I] @R1[I] @R1[P]
*#SAVE @C2[I] V(2) V(3) V(10) @R2[I] @R2[P] @RLOAD[I] @RLOAD[P]
*#SAVE V(5) V(4) @VIN[I] @VIN[P] V(6) @D2[ID] @D2[P]
*#ALIAS VSWITCHED  V(3)
*#VIEW  TRAN VSWITCHED
*#ALIAS VOUT  V(4)
*#VIEW  TRAN VOUT
.TRAN 100N 550U 500U 2N UIC
.OPTIONS ABSTOL=1U ITL1=1K METHOD=GEAR
.OPTIONS GMIN=100P RELTOL=0.005 VNTOL=1M
.OPTIONS MINSTEP=1N
.PRINT  TRAN VSWITCHED
.PRINT  TRAN VOUT
X2 2 6 FB 0 10 0 3 CS5171#0 
*{  }
.SUBCKT CS5171#0 VCC SYNC FB COM VC PGND VSW
*
X1 1 2 RAMP COM 5 3 X1_OSC#0 
*{  }
R9 5 16 100
X2 FB COM VC X2_ERRORAMP#0 
*{  }
R12 SYNC 19 500K
B1 3 COM V=1+TANH(1000*(V(VC)-V(SUM)))
R2 7 PGND 100K
R3 16 7 7
R4X 8 PGND 63M
Q3 VSW 7 8 Q2SC1847
.MODEL Q2SC1847 NPN BF=250 BR=4 CJC=82.8P CJE=256P IKF=.9
+ IKR=1.35 IS=152F ISE=60.8P MJC=.3 MJE=.5 NE=2 NF=1 NR=1
+ RB=.263 RC=26.3M RE=65.7M TF=1.06N TR=737N VAF=113 VAR=16
+ VJC=.3 VJE=1.1 XTB=1.5
B2 27 COM V=5*V(8)+.2*V(RAMP)+1.05
V2 19 COM DC=1.5
X4 VCC VCC COM 17 X_GATE#0 
*{  }
R4 22 20 100
B3 2 COM V=(56U+(2*56U)*(1+TANH(400*(V(FB)-.402))))*0.25*(V(ENABLE))
M1 23 20 COM COM SST211
.MODEL SST211 NMOS LEVEL=1 CBD=5.13E-12 CBS=6.16E-12
+ CGBO=2.34E-08 CGDO=3.00E-09 CGSO=3.60E-09 GAMMA=5.00E-06
+ IS=3.25E-14 KP=1.00E-02 LAMBDA=1.40E-02 MJ=.46 PB=0.80
+ PHI=0.75 RD=3.00E+01 RS=3.60E+01 TOX=3.00E-07 VTO=0.80
B4 22 COM V=1+TANH(100*(V(SYNC)-0.85))
C2 23 18 1N
X6 17 23 COM ENABLE X_GATE#0 
*{  }
R14 23 VCC 1MEG
B5 1 COM V=1+TANH(100*(V(SYNC)-2.5))
R11 23 18 100K
X8 17 17 COM 18 X_GATE#0 
*{  }
D3 16 VSW BAT83  M= 2
.MODEL BAT83 D BV=9.00E+01 CJO=1.31E-12 EG=0.69
+ IBV=1.00E-07 IS=9.98E-08 M=.333 N=1.47 RS=1.02E+01
+ TT=1.44E-11 VJ=.75 XTI=2
R16 SUM 27 1K
C4 SUM COM 10P
B7 VCC COM I=V(ENABLE) * (I(R3) * (1+0.002 * V(VCC)^2) + 0.25 * (6.2M + 0.023M 
+* V(VCC)))
B8 VCC COM I=25U * (8 + V(VCC)^2) / (40 + V(VCC)^2) - V(VCC) * 1U
.ENDS
C1 10 11 10NF
R1 11 0 5K
D2 3 4 1N5819
.MODEL 1N5819 D AF=1 BV=40 CJO=1.50114E-10 EG=1.3 FC=0.5
+ IBV=0.001 IS=1.19279E-05 KF=0 M=0.590203 N=1.16517
+ RS=0.0625421 TT=2.6273E-08 VJ=1.5 XTI=3.22098
C2 10 0 220PF
R2 2 6 1K
RLOAD 4 0 13
VIN 2 0 PULSE 0 3 0 100U
L2 2 1 22UH
R7 1 3 10M
R8 4 FB 3.72K
R9 FB 0 1.28K
C3 5 0 22UF
R10 4 5 100M
.SUBCKT X1_OSC#0 SYNC RATE RAMP COM Q R
C1 RAMP COM 100P
B1 3 COM V=TANH(100*(1-V(RAMP)+.5*V(2)))-.9
B2 COM RAMP I=V(RATE)*V(2)
R2 3 2 1
C2 2 COM 1N
X3 16 18 COM 13 X_GATE#0 
*{  }
B3 6 COM V=(1+TANH(1000*(.1-V(RAMP))))*2.5
R4 18 5 100
R3 RATE COM 1G
X4 R R COM 20 X_GATE#0 
*{  }
M1 RAMP 5 COM COM SST211
X5 13 6 COM 18 X_GATE#0 
*{  }
X6 SYNC 17 COM 16 X_GATE#0 
*{  }
X7 SYNC 4 COM 17 X_GATE#0 
*{  }
X1 9 Q COM 7 X_GATE#0 
*{  }
X2 7 12 COM Q X_GATE#0 
*{  }
R5 RAMP COM 10MEG
R6 6 9 1K
C3 9 COM 100P
X8 6 20 COM 12 X1_X8_GATE#0 
*{  }
R7 SYNC 4 1K
C5 4 COM 100P
.MODEL SST211 NMOS LEVEL=1 CBD=5.13E-12 CBS=6.16E-12
+ CGBO=2.34E-08 CGDO=3.00E-09 CGSO=3.60E-09 GAMMA=5.00E-06
+ IS=3.25E-14 KP=1.00E-02 LAMBDA=1.40E-02 MJ=.46 PB=0.80
+ PHI=0.75 RD=3.00E+01 RS=3.60E+01 TOX=3.00E-07 VTO=0.80
.MODEL Q2SC1847 NPN BF=250 BR=4 CJC=82.8P CJE=256P IKF=.9
+ IKR=1.35 IS=152F ISE=60.8P MJC=.3 MJE=.5 NE=2 NF=1 NR=1
+ RB=.263 RC=26.3M RE=65.7M TF=1.06N TR=737N VAF=113 VAR=16
+ VJC=.3 VJE=1.1 XTB=1.5
.MODEL SST211 NMOS LEVEL=1 CBD=5.13E-12 CBS=6.16E-12
+ CGBO=2.34E-08 CGDO=3.00E-09 CGSO=3.60E-09 GAMMA=5.00E-06
+ IS=3.25E-14 KP=1.00E-02 LAMBDA=1.40E-02 MJ=.46 PB=0.80
+ PHI=0.75 RD=3.00E+01 RS=3.60E+01 TOX=3.00E-07 VTO=0.80
.MODEL BAT83 D BV=9.00E+01 CJO=1.31E-12 EG=0.69
+ IBV=1.00E-07 IS=9.98E-08 M=.333 N=1.47 RS=1.02E+01
+ TT=1.44E-11 VJ=.75 XTI=2
.ENDS
.SUBCKT X2_ERRORAMP#0 FB COM OUT
B1 I1 COM V=SQRT((-25M-V(VFB))^2)*12
V5 7 0 DC=1.2
B3 COM OUT I=40U*TANH(SINH(V(I1))^1.5)-12U*V(I2)
B4 I2 COM V=EXPL(200*(5M+V(VFB)),1)
V3 VFB FB DC=-1.276
R1 FB COM 1G
D1 OUT 7 DN916
D2 7 OUT DN916
R3 OUT COM 1MEG
C1 OUT COM 120P
.MODEL DN916 D BV=133.3 CJO=1.75P IBV=10U IS=442P M=.333
+ N=1.70 RS=.42 TT=3.6N VJ=.75
.MODEL Q2SC1847 NPN BF=250 BR=4 CJC=82.8P CJE=256P IKF=.9
+ IKR=1.35 IS=152F ISE=60.8P MJC=.3 MJE=.5 NE=2 NF=1 NR=1
+ RB=.263 RC=26.3M RE=65.7M TF=1.06N TR=737N VAF=113 VAR=16
+ VJC=.3 VJE=1.1 XTB=1.5
.MODEL SST211 NMOS LEVEL=1 CBD=5.13E-12 CBS=6.16E-12
+ CGBO=2.34E-08 CGDO=3.00E-09 CGSO=3.60E-09 GAMMA=5.00E-06
+ IS=3.25E-14 KP=1.00E-02 LAMBDA=1.40E-02 MJ=.46 PB=0.80
+ PHI=0.75 RD=3.00E+01 RS=3.60E+01 TOX=3.00E-07 VTO=0.80
.MODEL BAT83 D BV=9.00E+01 CJO=1.31E-12 EG=0.69
+ IBV=1.00E-07 IS=9.98E-08 M=.333 N=1.47 RS=1.02E+01
+ TT=1.44E-11 VJ=.75 XTI=2
.ENDS
.SUBCKT X_GATE#0 A B COM OUT
R1 A B 1MEG
B1 3 COM V=(1+TANH(1000*(1.5-V(A))))*(1+TANH(1000*(1.5-V(B))))
R2 3 OUT 1
C1 OUT COM 1N
.MODEL Q2SC1847 NPN BF=250 BR=4 CJC=82.8P CJE=256P IKF=.9
+ IKR=1.35 IS=152F ISE=60.8P MJC=.3 MJE=.5 NE=2 NF=1 NR=1
+ RB=.263 RC=26.3M RE=65.7M TF=1.06N TR=737N VAF=113 VAR=16
+ VJC=.3 VJE=1.1 XTB=1.5
.MODEL SST211 NMOS LEVEL=1 CBD=5.13E-12 CBS=6.16E-12
+ CGBO=2.34E-08 CGDO=3.00E-09 CGSO=3.60E-09 GAMMA=5.00E-06
+ IS=3.25E-14 KP=1.00E-02 LAMBDA=1.40E-02 MJ=.46 PB=0.80
+ PHI=0.75 RD=3.00E+01 RS=3.60E+01 TOX=3.00E-07 VTO=0.80
.MODEL BAT83 D BV=9.00E+01 CJO=1.31E-12 EG=0.69
+ IBV=1.00E-07 IS=9.98E-08 M=.333 N=1.47 RS=1.02E+01
+ TT=1.44E-11 VJ=.75 XTI=2
.ENDS
.SUBCKT X1_X8_GATE#0 A B COM OUT
R1 A B 1MEG
B1 3 COM V=4-(1+TANH(1000*(1.5-V(A))))*(1+TANH(1000*(1.5-V(B))))
R2 3 OUT 1
C1 OUT COM 1N
.MODEL Q2SC1847 NPN BF=250 BR=4 CJC=82.8P CJE=256P IKF=.9
+ IKR=1.35 IS=152F ISE=60.8P MJC=.3 MJE=.5 NE=2 NF=1 NR=1
+ RB=.263 RC=26.3M RE=65.7M TF=1.06N TR=737N VAF=113 VAR=16
+ VJC=.3 VJE=1.1 XTB=1.5
.MODEL SST211 NMOS LEVEL=1 CBD=5.13E-12 CBS=6.16E-12
+ CGBO=2.34E-08 CGDO=3.00E-09 CGSO=3.60E-09 GAMMA=5.00E-06
+ IS=3.25E-14 KP=1.00E-02 LAMBDA=1.40E-02 MJ=.46 PB=0.80
+ PHI=0.75 RD=3.00E+01 RS=3.60E+01 TOX=3.00E-07 VTO=0.80
.MODEL BAT83 D BV=9.00E+01 CJO=1.31E-12 EG=0.69
+ IBV=1.00E-07 IS=9.98E-08 M=.333 N=1.47 RS=1.02E+01
+ TT=1.44E-11 VJ=.75 XTI=2
.ENDS
.END
